// 115200 bits per second = 8.68us
`define BAUD 115200
// 25MHz = 40ns period
`define SOURCE_FREQ 25000000
// Bit size of accumulator
`define ACCUMULATOR_WIDTH 16

// Uncomment if you want to use 1 stop bit
`define ONE_STOP_BIT
// `define TWO_STOP_BITS
