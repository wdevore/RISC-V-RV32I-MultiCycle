`define MEM_WORDS 4
`define DATA_WIDTH 8
