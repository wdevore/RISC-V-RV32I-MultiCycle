
typedef enum logic [3:0] {
    Idle,
    Transmitting,
    Complete,
    Reset
} TxState /*verilator public*/; 
