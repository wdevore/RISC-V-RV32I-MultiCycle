
typedef enum logic [3:0] {
    CSReset,
    CSReset1,
    CSResetComplete
} ControlState; 

