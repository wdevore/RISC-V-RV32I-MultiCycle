`define RESET_VECTOR 32'h00000300

// For embedded memory contents
`define ROM_PATH "../rams/"
`define MEM_CONTENTS "code"
`define ROM_EXTENSION ".ram"
